PACKAGE harq_type IS

    TYPE HARQ_RESP IS(ACK_T1, ACK_T2, NACK);

END PACKAGE harq_type;