PACKAGE harq_type IS

    TYPE HARQ_RESP IS(ACK, NACK);

END PACKAGE harq_type;