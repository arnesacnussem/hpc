PACKAGE decoder_types IS
    TYPE DecoderType IS (PMS2, BAO3, UNDEFINED);
END PACKAGE decoder_types;