
LIBRARY ieee;
PACKAGE consts IS
    CONSTANT MSG_LENGTH : INTEGER := 10; --	msg len = 11
    CONSTANT CODEWORD_LENGTH : INTEGER := 14; --	codeword len = 15
    CONSTANT CHK_LENGTH : INTEGER := 3; --	check bits = 4
    TYPE GEN_MAT IS ARRAY (0 TO MSG_LENGTH, 0 TO CODEWORD_LENGTH) OF BIT;
    TYPE CHK_MAT IS ARRAY (0 TO CHK_LENGTH, 0 TO CODEWORD_LENGTH) OF BIT;
    TYPE MSG_ENC IS ARRAY(0 TO CODEWORD_LENGTH) OF BIT;
    TYPE MESSAGE IS ARRAY (0 TO MSG_LENGTH) OF BIT;
    CONSTANT GENERATE_MATRIX : GEN_MAT := (
        0 => "110010000000000",
		1 => "011001000000000",
		2 => "001100100000000",
		3 => "110100010000000",
		4 => "101000001000000",
		5 => "010100000100000",
		6 => "111000000010000",
		7 => "011100000001000",
		8 => "111100000000100",
		9 => "101100000000010",
		10 => "100100000000001"
    );
    CONSTANT CHECK_MATRIX : CHK_MAT := (
        0 => "100010011010111",
		1 => "010011010111100",
		2 => "001001101011110",
		3 => "000100110101111"
    );
END PACKAGE consts;
