LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
PACKAGE consts IS
    CONSTANT MSG_LENGTH : INTEGER := 4 - 1;
    CONSTANT CODEWORD_LENGTH : INTEGER := 7 - 1;
    TYPE GEN_MAT IS ARRAY (0 TO MSG_LENGTH, 0 TO CODEWORD_LENGTH) OF BIT;
    TYPE CHK_MAT IS ARRAY (0 TO MSG_LENGTH, 0 TO CODEWORD_LENGTH) OF BIT;
    TYPE MSG_ENC IS ARRAY(0 TO CODEWORD_LENGTH) OF BIT;
    TYPE MESSAGE IS ARRAY (0 TO MSG_LENGTH) OF BIT;
END PACKAGE consts;