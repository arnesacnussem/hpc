LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY trransport IS
    PORT (
        clk, en : IN STD_LOGIC;
        dat_in  : IN BIT;
        dat_out : OUT BIT
    );
END trransport;

ARCHITECTURE Transportor OF trransport IS

BEGIN
 
END ARCHITECTURE;