
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
PACKAGE consts IS
    CONSTANT MSG_LENGTH : INTEGER := 3; --	msg len = 4
    CONSTANT CODEWORD_LENGTH : INTEGER := 6; --	codeword len = 7
    CONSTANT CHK_LENGTH : INTEGER := 2; --	check bits = 3
    TYPE GEN_MAT IS ARRAY (0 TO MSG_LENGTH, 0 TO CODEWORD_LENGTH) OF BIT;
    TYPE CHK_MAT IS ARRAY (0 TO CHK_LENGTH, 0 TO CODEWORD_LENGTH) OF BIT;
    TYPE MSG_ENC IS ARRAY(0 TO CODEWORD_LENGTH) OF BIT;
    TYPE MESSAGE IS ARRAY (0 TO MSG_LENGTH) OF BIT;
    CONSTANT GENERATE_MATRIX : GEN_MAT := (
        0 => "1101000",
		1 => "0110100",
		2 => "1110010",
		3 => "1010001"
    );
    CONSTANT CHECK_MATRIX : CHK_MAT := (
        0 => "1001011",
		1 => "0101110",
		2 => "0010111"
    );
END PACKAGE consts;
