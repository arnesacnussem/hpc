PACKAGE decoder_types IS
    TYPE DecoderType IS (PMS2, BAO3, DUMMY);
END PACKAGE decoder_types;