LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
PACKAGE consts IS
    CONSTANT MSG_LENGTH : INTEGER := 4 - 1;
    CONSTANT CODEWORD_LENGTH : INTEGER := 7 - 1;
    TYPE generator_matrix IS ARRAY (0 TO MSG_LENGTH, 0 TO CODEWORD_LENGTH) OF BIT;
    TYPE code_matrix IS ARRAY (0 TO CODEWORD_LENGTH, 0 TO MSG_LENGTH) OF BIT;
    TYPE code_matrix_transpose IS ARRAY (0 TO MSG_LENGTH, 0 TO CODEWORD_LENGTH) OF BIT;
END PACKAGE consts;