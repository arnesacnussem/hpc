PACKAGE consts IS
    CONSTANT MSG_LENGTH : INTEGER := 4 - 1;
    CONSTANT CODEWORD_LENGTH : INTEGER := 7 - 1;
    TYPE generator_matrix IS ARRAY (CODEWORD_LENGTH DOWNTO 0, MSG_LENGTH DOWNTO 0) OF BIT;
    TYPE code_matrix IS ARRAY (CODEWORD_LENGTH DOWNTO 0, MSG_LENGTH DOWNTO 0) OF BIT;
    TYPE code_matrix_transpose IS ARRAY (MSG_LENGTH DOWNTO 0, CODEWORD_LENGTH DOWNTO 0) OF BIT;
END PACKAGE consts;