LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.math_real.ALL;
USE work.generated.ALL;

ENTITY encoder_mxio IS
    GENERIC (
        MSG_RATIO  : POSITIVE := MSG_SERIAL'length;
        CODE_RATIO : POSITIVE := CODEWORD_SERIAL'length;
        -- [0]: 输入缓存
        -- [1]: 输出填充
        IO_CONTROL : BIT_VECTOR(0 TO 1) := "10"
    );
    PORT (
        msg   : IN BIT_VECTOR(0 TO MSG_SERIAL'length / MSG_RATIO - 1);
        code  : OUT BIT_VECTOR(0 TO CODEWORD_SERIAL'length / CODE_RATIO - 1);
        clk   : IN STD_LOGIC;
        ready : OUT STD_LOGIC
    );
END ENTITY;

ARCHITECTURE encoder_mxio OF encoder_mxio IS
    SIGNAL msg_matrix  : MSG_MAT;
    SIGNAL code_matrix : CODEWORD_MAT;
    SIGNAL rst         : STD_LOGIC              := '0';
    SIGNAL in_port     : BIT_VECTOR(msg'RANGE)  := msg;
    SIGNAL out_port    : BIT_VECTOR(code'RANGE) := code;

    -- [0] mxio_in_ready
    -- [1] codec_ready
    -- [2] mxio_out_ready
    SIGNAL state : STD_ULOGIC_VECTOR(0 TO 2) := "000";

    -- clock control
    SIGNAL mxio_in_clk  : STD_LOGIC;
    SIGNAL codec_clk    : STD_LOGIC;
    SIGNAL mxio_out_clk : STD_LOGIC;

BEGIN
    enc_mxio_in : ENTITY work.matrix_io
        GENERIC MAP(
            COL_CNT  => MSG_LINE'length,
            ROW_CNT  => MSG_MAT'length,
            IO_WIDTH => msg'length,
            IO_MODE  => '0' & IO_CONTROL(0)
        )
        PORT MAP(
            io_port => in_port,
            matrix  => msg_matrix,
            clk     => mxio_in_clk,
            ready   => state(0)
        );

    encoder_inst : ENTITY work.encoder
        PORT MAP(
            msg   => msg_matrix,
            code  => code_matrix,
            ready => state(1),
            rst   => rst,
            clk   => codec_clk
        );
    enc_mxio_out : ENTITY work.matrix_io
        GENERIC MAP(
            COL_CNT  => CODEWORD_LINE'length,
            ROW_CNT  => CODEWORD_MAT'length,
            IO_WIDTH => code'length,
            IO_MODE  => '1' & IO_CONTROL(1)
        )
        PORT MAP(
            io_port => out_port,
            matrix  => code_matrix,
            clk     => mxio_out_clk,
            ready   => state(2)
        );
    PROCESS (ALL)
    BEGIN
        in_port <= msg;
        code    <= out_port;
        ready   <= state(2);
        CASE state IS
            WHEN "000" =>
                mxio_in_clk  <= clk;
                codec_clk    <= '0';
                mxio_out_clk <= '0';
            WHEN "100" =>
                mxio_in_clk  <= '0';
                codec_clk    <= clk;
                mxio_out_clk <= '0';
            WHEN "110" =>
                mxio_in_clk  <= '0';
                codec_clk    <= '0';
                mxio_out_clk <= clk;
            WHEN OTHERS =>
                mxio_in_clk  <= '0';
                codec_clk    <= '0';
                mxio_out_clk <= '0';
        END CASE;
    END PROCESS;

END ARCHITECTURE;