PACKAGE decoder_types IS
    TYPE DecoderType IS (EHPC, SHPC, BAO3, DUMMY);
END PACKAGE decoder_types;